LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY register8 IS
	PORT(
		Clock:IN STD_LOGIC;
		RESET:IN STD_LOGIC ;
		INPUT:IN STD_LOGIC_VECTOR(0 TO 7);
		OUTPUT:OUT STD_LOGIC_VECTOR(0 TO 7) 
	);
END register8;

ARCHITECTURE content OF register8 IS

BEGIN
	PROCESS(RESET , Clock) --sensitive signal
	BEGIN 
	
	IF  RESET = '0' THEN 
		OUTPUT <= "00000000";
	ELSIF rising_edge (Clock) THEN
		OUTPUT <= INPUT;
	END IF;
	END PROCESS;
	
END content;