LIBRARY ieee;
USE ieee.std_logic_1164.all;


ENTITY  trans416 IS
	PORT
	(
		A:IN STD_LOGIC_VECTOR(3 downto 0);
		EN: IN STD_LOGIC;
		Y: OUT STD_LOGIC_VECTOR(15 downto 0)
	);
END trans416;

ARCHITECTURE dec_behave OF  trans416 IS
signal sel: STD_LOGIC_VECTOR(4 downto 0);

BEGIN
	sel <= A&EN;
	WITH sel SELECT
	Y<= "1111111111111110" WHEN "00001",
		"1111111111111101" WHEN "00011",
		"1111111111111011" WHEN "00101",
		"1111111111110111" WHEN "00111",
		"1111111111101111" WHEN "01001",
		"1111111111011111" WHEN "01011",
		"1111111110111111" WHEN "01101",
		"1111111101111111" WHEN "01111",
		"1111111011111111" WHEN "10001",
		"1111110111111111" WHEN "10011",
		"1111101111111111" WHEN "10101",
		"1111011111111111" WHEN "10111",
		"1110111111111111" WHEN "11001",
		"1101111111111111" WHEN "11011",
		"1011111111111111" WHEN "11101",
		"0111111111111111" WHEN "11111",
		"1111111111111111" WHEN OTHERS;		
END  dec_behave;
