LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY encode83 IS
	PORT(
		D:IN STD_LOGIC_VECTOR(0 TO 7);
		A:OUT STD_LOGIC_VECTOR(0 TO 2)
	);
END encode83;

ARCHITECTURE content OF encode83 IS
BEGIN
PROCESS(D)
BEGIN 
 IF	(D(7)='0') THEN A<="111";
	ELSIF (D(6)='0') THEN A<="110";
	ELSIF (D(5)='0') THEN A<="101";
	ELSIF (D(4)='0') THEN A<="100";
	ELSIF (D(3)='0') THEN A<="011";
	ELSIF (D(2)='0') THEN A<="010";
	ELSIF (D(1)='0') THEN A<="001";
	ELSIF (D(0)='0') THEN A<="000";
	ELSE A<="ZZZ";
	END IF;
END PROCESS;
END;